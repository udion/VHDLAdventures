----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:05:17 01/30/2017 
-- Design Name: 
-- Module Name:    encrypter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity encrypter is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           plaintext : in  STD_LOGIC_VECTOR (63 downto 0);
           start : in  STD_LOGIC;
           ciphertext : out  STD_LOGIC_VECTOR (63 downto 0);
           done : out  STD_LOGIC);
end encrypter;

architecture Behavioral of encrypter is
constant key:STD_LOGIC_VECTOR (127 downto 0) := x"ff0f745743fd99f775f8c48f2927c18c";
constant k0: STD_LOGIC_VECTOR (31 downto 0):= key(31 downto 0);
constant k1: STD_LOGIC_VECTOR (31 downto 0) := key(63 downto 32);
constant k2: STD_LOGIC_VECTOR (31 downto 0) := key(95 downto 64);
constant k3: STD_LOGIC_VECTOR (31 downto 0) := key(127 downto 96);
constant delta : STD_LOGIC_VECTOR (31 downto 0):=x"9E3779B9";

signal sum: STD_LOGIC_VECTOR (31 downto 0):=x"00000000";
signal cv0,cv1: std_logic_vector (31 downto 0);
signal temp1,temp2,temp3,temp4:STD_LOGIC_VECTOR (31 downto 0):= (others => '0');
signal counter :integer:=0;
begin
	process(clk, start,reset)
	begin
		if(reset='1') then
			ciphertext<=(others=>'0');
			done<='0';
		else
			if (clk='1') then
					if (start='1') then
						if(counter = 0) then
							cv0 <= plaintext(31 downto 0);
							cv1 <= plaintext(63 downto 32);
							done <= '0';
						elsif (counter<97 and (counter mod 3 = 1)) then
							sum <= sum+delta;
						elsif (counter<97 and (counter mod 3 = 2)) then
							cv0 <= cv0+(((cv1(27 downto 0) & "0000")+k0)xor(cv1+sum)xor(("00000" & cv1(31 downto 5))+k1));
						elsif (counter<97 and (counter mod 3 = 0)) then
							cv1 <= cv1+(((cv0(27 downto 0) & "0000")+k2)xor(cv0+sum)xor(("00000" & cv0(31 downto 5))+k3));
						else
							ciphertext <= cv1&cv0;
							done<='1';
						end if;
					counter <= counter+1;
					end if;
			end if;
		end if;
	end process;
end Behavioral;